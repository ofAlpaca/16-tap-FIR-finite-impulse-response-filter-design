module rom(out, cs, address, clk);
	input cs, clk;
	input [4:0]address;
	output [7:0]out;
	
	reg [7:0]out;
	reg [7:0]a[0:31];
	/*
	always@(posedge clk) begin
			case(address)
				5'd0: c[0] = 8'b0_1000000;
				5'd1: c[1] = 8'b0_0100000;
				5'd2: c[2] = 8'b0_1100000;
				5'd3: c[3] = 8'b0_0010000;
				5'd4: c[4] = 8'b0_1010000;
				5'd5: c[5] = 8'b0_0110000;
				5'd6: c[6] = 8'b0_1110000;
				5'd7: c[7] = 8'b0_0001000;
				5'd8: c[8] = 8'b0_1001000;
				5'd9: c[9] = 8'b0_0101000;
				5'd10: c[10] = 8'b0_1101000;
				5'd11: c[11] = 8'b0_0011000;
				5'd12: c[12] = 8'b0_1011000;
				5'd13: c[13] = 8'b0_0111000;
				5'd14: c[14] = 8'b0_1111000;
				5'd15: c[15] = 8'b0_0000100;
				5'd31: c[31] = 8'b1_0000000;
				default: c[address] = 0;
			endcase
		
	end
	
	assign out = cs? c[address]:8'hxx;
	*/
	always@(posedge clk) begin
			case(address)
				5'd0: a[0] = 8'b0_1110011;
				5'd1: a[1] = 8'b0_0110100;
				5'd2: a[2] = 8'b0_1110100;
				5'd3: a[3] = 8'b0_0011001;
				5'd4: a[4] = 8'b0_1010111;
				5'd5: a[5] = 8'b1_1110001;
				5'd6: a[6] = 8'b0_1010110;
				5'd7: a[7] = 8'b0_0000100;
				5'd8: a[8] = 8'b1_0000101;
				5'd9: a[9] = 8'b1_1100000;
				5'd10: a[10] = 8'b0_1100110;
				5'd11: a[11] = 8'b1_1101101;
				5'd12: a[12] = 8'b1_0110011;
				5'd13: a[13] = 8'b1_1001101;
				5'd14: a[14] = 8'b0_0001001;
				5'd15: a[15] = 8'b0_1101001;
				5'd16: a[16] = 8'b0_0000110;
				5'd17: a[17] = 8'b1_1001110;
				5'd18: a[18] = 8'b1_0001000;
				5'd19: a[19] = 8'b0_0110111;
				5'd20: a[20] = 8'b0_1000100;
				5'd21: a[21] = 8'b1_0001111;
				5'd22: a[22] = 8'b0_0100000;
				5'd23: a[23] = 8'b1_1000011;
				5'd24: a[24] = 8'b1_1001111;
				5'd25: a[25] = 8'b0_0000101;
				5'd26: a[26] = 8'b1_1101000;
				5'd27: a[27] = 8'b0_1100100;
				5'd28: a[28] = 8'b0_0010010;
				5'd29: a[29] = 8'b0_0010001;
				5'd30: a[30] = 8'b1_1100100;
				5'd31: a[31] = 8'b0_0110001;
			endcase
		
		if(cs)
			out = a[address];
		else
			out = 8'bxxxxxxxx;
	end
endmodule